module main

fn grains_on_square(square int) !u64 {
}

fn total_grains_on_board() u64 {
	// totally unnessesary comment
}
